library ieee;
use ieee.std_logic_1164.all;

package start_condition_graphic is
    constant start_condition_width : integer := 299;
    constant start_condition_height : integer := 15;
    type start_condition_array is array (0 to start_condition_height-1, 0 to start_condition_width-1) of std_logic_vector(11 downto 0);
    constant START_CONDITION_IMAGE : start_condition_array := (
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"EEE", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"EEE", X"EEE", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"EEE", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"EEE", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"EEE", X"EEE", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"EEE", X"EEE", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"FFF", X"EEE", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"EEE", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"EEE", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"EEE", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"DDD", X"EEE", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"EEE", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"DDD", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"111", X"444", X"444", X"444", X"111", X"000", X"000", X"222", X"FFF", X"BBB", X"000", X"000", X"000", X"333", X"444", X"444", X"333", X"000", X"000", X"000", X"555", X"FFF", X"666", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"444", X"444", X"CCC", X"FFF", X"222", X"000", X"000", X"111", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"FFF", X"BBB", X"000", X"000", X"000", X"222", X"444", X"444", X"444", X"444", X"444", X"333", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"111", X"444", X"444", X"444", X"444", X"444", X"444", X"666", X"FFF", X"999", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"444", X"333", X"AAA", X"FFF", X"888", X"333", X"444", X"444", X"000", X"000", X"000", X"111", X"444", X"444", X"444", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"333", X"444", X"444", X"333", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"333", X"444", X"444", X"222", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"333", X"444", X"444", X"333", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"222", X"444", X"444", X"444", X"333", X"666", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"666", X"333", X"444", X"333", X"000", X"000", X"000", X"222", X"444", X"444", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"333", X"444", X"444", X"000", X"000", X"000", X"111", X"444", X"444", X"333", X"BBB", X"FFF", X"222", X"000", X"000", X"111", X"444", X"444", X"444", X"111", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"444", X"333", X"BBB", X"FFF", X"666", X"333", X"444", X"333", X"000", X"000", X"000", X"222", X"444", X"444", X"444", X"FFF", X"DDD", X"000", X"000", X"000", X"222", X"444", X"444", X"444", X"000", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"333", X"444", X"444", X"333", X"000", X"000", X"000", X"999", X"FFF", X"777", X"333", X"444", X"333", X"000", X"000", X"000", X"222", X"444", X"444", X"444"),
    (X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"222", X"FFF", X"BBB", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"444", X"BBB", X"AAA", X"BBB", X"333", X"000", X"000", X"222", X"FFF", X"BBB", X"000", X"000", X"000", X"777", X"BBB", X"BBB", X"AAA", X"000", X"000", X"000", X"666", X"FFF", X"666", X"000", X"000", X"000", X"AAA", X"BBB", X"AAA", X"BBB", X"AAA", X"DDD", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"333", X"BBB", X"AAA", X"AAA", X"AAA", X"BBB", X"EEE", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"666", X"BBB", X"AAA", X"BBB", X"AAA", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"444", X"BBB", X"AAA", X"AAA", X"AAA", X"BBB", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"777", X"BBB", X"AAA", X"BBB", X"AAA", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"AAA", X"AAA", X"BBB", X"666", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"777", X"BBB", X"BBB", X"999", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"CCC", X"AAA", X"BBB", X"BBB", X"AAA", X"CCC", X"FFF", X"777", X"000", X"000", X"000", X"999", X"BBB", X"BBB", X"777", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"999", X"BBB", X"AAA", X"BBB", X"AAA", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"999", X"BBB", X"BBB", X"777", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"333", X"000", X"000", X"000", X"000", X"555", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"999", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"777", X"AAA", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"999", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"888", X"FFF", X"DDD", X"888", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"777", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"888", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"777", X"BBB", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"444", X"000", X"000", X"000", X"000", X"666", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"777", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"888", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"333", X"888", X"777", X"777", X"111", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"777", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"333", X"000", X"000", X"000", X"000", X"555", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"333", X"999", X"888", X"999", X"888", X"999", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"666", X"999", X"999", X"888", X"000", X"111", X"666", X"AAA", X"FFF", X"666", X"000", X"000", X"000", X"888", X"999", X"888", X"999", X"888", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"999", X"888", X"888", X"888", X"999", X"333", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"DDD", X"888", X"888", X"888", X"999", X"888", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"333", X"999", X"888", X"888", X"888", X"999", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"666", X"999", X"888", X"999", X"888", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"888", X"999", X"999", X"555", X"000", X"444", X"777", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"666", X"999", X"999", X"777", X"000", X"111", X"666", X"BBB", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"AAA", X"888", X"000", X"000", X"000", X"555", X"FFF", X"777", X"000", X"000", X"000", X"777", X"999", X"999", X"666", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"888", X"999", X"888", X"999", X"666", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"777", X"999", X"999", X"666", X"000", X"222", X"666", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"555", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"555", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"666", X"FFF", X"666", X"000", X"000", X"000", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"CCC", X"FFF", X"666", X"444", X"444", X"444", X"444", X"444", X"444", X"111", X"000", X"000", X"000", X"FFF", X"CCC", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"111", X"444", X"444", X"444", X"444", X"444", X"EEE", X"FFF", X"000", X"000", X"000", X"111", X"444", X"444", X"444", X"444", X"444", X"444", X"666", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"333", X"444", X"444", X"333", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"EEE", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"222", X"444", X"444", X"333", X"000", X"000", X"000", X"555", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"111", X"444", X"444", X"444", X"111", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"333", X"444", X"444", X"444", X"444", X"444", X"333", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"555", X"CCC", X"BBB", X"BBB", X"111", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"CCC", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"BBB", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"DDD", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"CCC", X"DDD", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"EEE", X"DDD", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"BBB", X"DDD", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"DDD", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"555", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"444", X"FFF", X"777", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF")
    );
end package start_condition_graphic;
