library ieee;
use ieee.std_logic_1164.all;

package brown_car_image_graphic is
    constant BROWN_CAR_IMAGE : array (0 to 87, 0 to 65) of std_logic_vector(11 downto 0) := (
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FD3", X"FD3", X"FD3", X"FD3", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FD3", X"FD3", X"FD3", X"FD3", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FD3", X"FD3", X"FD3", X"FD3", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FD3", X"FD3", X"FD3", X"FD3", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FD3", X"FD3", X"FD3", X"FD3", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FD3", X"FD3", X"FD3", X"FD3", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FD3", X"FD3", X"FD3", X"FD3", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FD3", X"FD3", X"FD3", X"FD3", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"832", X"832", X"832", X"832", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"A53", X"A53", X"A53", X"A53", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"FD3", X"FD3", X"FD3", X"FD3", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"074", X"A53", X"A53", X"A53", X"A53", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    );
end package;
