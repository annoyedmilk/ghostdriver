library ieee;
use ieee.std_logic_1164.all;

package game_over_graphic is
    constant game_over_width : integer := 305;
    constant game_over_height : integer := 42;
    type game_over_array is array (0 to game_over_height-1, 0 to game_over_width-1) of std_logic_vector(11 downto 0);
    constant GAME_OVER_IMAGE : game_over_array := (
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"333", X"333", X"333", X"333", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"333", X"333", X"333", X"333", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"777", X"777", X"777", X"777", X"777", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"888", X"777", X"777", X"777", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"777", X"777", X"888", X"777", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"111", X"777", X"777", X"777", X"777", X"777", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"888", X"777", X"888", X"777", X"777", X"111", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"777", X"888", X"777", X"777", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"777", X"777", X"888", X"777", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"777", X"777", X"777", X"777", X"777"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"BBB", X"BBB", X"BBB", X"BBB", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"BBB", X"BBB", X"BBB", X"BBB", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"EEE", X"EEE", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"777", X"777", X"777", X"777", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"777", X"777", X"777", X"777", X"333", X"000", X"000", X"000", X"000", X"222", X"777", X"777", X"777", X"777", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"888", X"777", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"888", X"777", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"333", X"000", X"000", X"000", X"000", X"222", X"777", X"777", X"777", X"777", X"777"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"444", X"444", X"444", X"444", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"AAA", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"444", X"444", X"444", X"444", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000")
    );
end package game_over_graphic;
