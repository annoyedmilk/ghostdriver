library ieee;
use ieee.std_logic_1164.all;

package blue_car_graphic is
		constant blue_car_width : integer := 66;
    constant blue_car_height : integer := 88;
    type blue_car_array is array (0 to blue_car_height-1, 0 to blue_car_width-1) of std_logic_vector(11 downto 0);
    constant BLUE_CAR_IMAGE : blue_car_array := (
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"074", X"074", X"074", X"074", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"074", X"074", X"074", X"074", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"074", X"074", X"074", X"074", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"074", X"074", X"074", X"074", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"074", X"074", X"074", X"074", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"074", X"074", X"074", X"074", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"074", X"074", X"074", X"074", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"074", X"074", X"074", X"074", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"4AC", X"4AC", X"4AC", X"4AC", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"23D", X"4AC", X"4AC", X"4AC", X"4AC", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
        (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB")
    );
end package blue_car_graphic;
