library ieee;
use ieee.std_logic_1164.all;

package ghost_driver_graphic is
    constant ghost_driver_width : integer := 389;
    constant ghost_driver_height : integer := 42;
    type ghost_driver_array is array (0 to ghost_driver_height-1, 0 to ghost_driver_width-1) of std_logic_vector(11 downto 0);
    constant GHOST_DRIVER_IMAGE : ghost_driver_array := (
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"444", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"333", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"777", X"777", X"777", X"777", X"777", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"777", X"888", X"777", X"777", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"777", X"777", X"777", X"777", X"777", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"777", X"888", X"777", X"777", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"777", X"777", X"888", X"777", X"888", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"777", X"777", X"888", X"777", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"777", X"777", X"777", X"777", X"777"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"444", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"BBB", X"BBB", X"BBB", X"BBB", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"444", X"444", X"444", X"444", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"BBB", X"BBB", X"BBB", X"BBB", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"777", X"777", X"777", X"777", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"777", X"888", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"222", X"000", X"000", X"000", X"000", X"333", X"777", X"777", X"888", X"777", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"888", X"777", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"777", X"333", X"000", X"000", X"000", X"000", X"222", X"777", X"777", X"777", X"777", X"777"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"888", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"888", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"DDD", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"AAA", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"444", X"444", X"444", X"444", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"444", X"444", X"444", X"444", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"999", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"000", X"777", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"999", X"000", X"111", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"DDD", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"333", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"444", X"FFF", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"EEE", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"EEE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
    (X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"AAA", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"CCC", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"555", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"444", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"333", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"555", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"222", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"222", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"666", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"666", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"AAA", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"CCC", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"111", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"777", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000")
    );
end package ghost_driver_graphic;
