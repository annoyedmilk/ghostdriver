constant BLACK_CAR_IMAGE : array (0 to 87, 0 to 65) of std_logic_vector(11 downto 0) := (
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"E86", X"E86", X"E86", X"E86", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"E86", X"E86", X"E86", X"E86", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"E86", X"E86", X"E86", X"E86", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"E86", X"E86", X"E86", X"E86", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"E86", X"E86", X"E86", X"E86", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"E86", X"E86", X"E86", X"E86", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"E86", X"E86", X"E86", X"E86", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"E86", X"E86", X"E86", X"E86", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
);
