library ieee;
use ieee.std_logic_1164.all;

package black_car_graphic is
    constant car_width : integer := 66;
    constant car_height : integer := 88;
    type black_car_array is array (0 to car_height-1, 0 to car_width-1) of std_logic_vector(11 downto 0);
    constant BLACK_CAR_IMAGE : black_car_array := (
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"000", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"000", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"000", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"000", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"E86", X"E86", X"E86", X"E86", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"E86", X"E86", X"E86", X"E86", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"E86", X"E86", X"E86", X"E86", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"E86", X"E86", X"E86", X"E86", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FFF", X"FFF", X"FFF", X"FFF", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"527", X"527", X"527", X"527", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"527", X"527", X"527", X"527", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB")
    );
end package black_car_graphic;
