constant RED_CAR_IMAGE : array (0 to 87, 0 to 65) of std_logic_vector(11 downto 0) := (
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E86", X"E86", X"E86", X"E86", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"566", X"566", X"566", X"566", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"566", X"566", X"566", X"566", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"566", X"566", X"566", X"566", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"566", X"566", X"566", X"566", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"566", X"566", X"566", X"566", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"566", X"566", X"566", X"566", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"566", X"566", X"566", X"566", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"566", X"566", X"566", X"566", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"832", X"E86", X"E86", X"E86", X"E86", X"000", X"000", X"000", X"000", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E86", X"E36", X"E36", X"E36", X"E36", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"832", X"832", X"832", X"832", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"FD3", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"E36", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"566", X"566", X"566", X"566", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"566", X"A53", X"A53", X"A53", X"A53", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
    (X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB", X"BBB"),
);
